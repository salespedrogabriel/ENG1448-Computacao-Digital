use IEEE.STD_LOGIC_1164.ALL;

entity u_estados is
end u_estados;

architecture Behavioral of u_estados is

begin


end Behavioral;

